module Adder16bit(input[15:0] A, B, output[15:0] W);
	wire[15:0] c;
	FA f1(A[0], B[0], 1'b0, W[0], c[0]);
	FA f2(A[1], B[1], c[0], W[1], c[1]);
	FA f3(A[2], B[2], c[1], W[2], c[2]);
	FA f4(A[3], B[3], c[2], W[3], c[3]);
	FA f5(A[4], B[4], c[3], W[4], c[4]);
	FA f6(A[5], B[5], c[4], W[5], c[5]);
	FA f7(A[6], B[6], c[5], W[6], c[6]);
	FA f8(A[7], B[7], c[6], W[7], c[7]);
	FA f9(A[8], B[8], c[7], W[8], c[8]);
	FA f10(A[9], B[9], c[8], W[9], c[9]);
	FA f11(A[10], B[10], c[9], W[10], c[10]);
	FA f12(A[11], B[11], c[10], W[11], c[11]);
	FA f13(A[12], B[12], c[11], W[12], c[12]);
	FA f14(A[13], B[13], c[12], W[13], c[13]);
	FA f15(A[14], B[14], c[13], W[14], c[14]);
	FA f16(A[15], B[15], c[14], W[15], c[15]);
endmodule
